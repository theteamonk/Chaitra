/********************************************************************************************
Filename    :	    router_fifo.v   

Description :      FIFO 16x9 sublock Design

Author Name :      Chaitra

Version     :      1.0

Width allocation:
  8     7 6 5 4 3 2    1 0
parity    payload     header
********************************************************************************************/

module router_fifo(clock, resetn, data_in, read_enb, write_enb, 
			data_out, full, empty, lfd_state, soft_reset);

parameter width = 9,
	  depth = 16;
	  
input lfd_state;
input [width-2 : 0] data_in;
input clock, resetn, read_enb, write_enb, soft_reset;

output reg [width-2 : 0] data_out;
output full, empty;

reg [4:0] rd_ptr, wr_ptr;		//internal pointers
reg [6:0] count;			//internal counter
reg [width-1 : 0] mem [depth-1 : 0];	//memory declaration
reg temp;				//to delay the lfd_state bit by one clock cycle

integer i;

/******************************************fifo full and empty logic**************************************************/
/*???check if full and empty logic can be written in a different way???*/

//combinational logic
//empty flag
//when write pointer and read pointer are pointing at the same location, empty = 1. Continuous check is needed
assign empty = (wr_ptr == rd_ptr);	

//full flag
//when the locations are filled with data and write pointer increments to the 16th location (as it is a 5-bit pointer)
//and read pointer still not started to point and read the data (still in 0th location)
//vector slicing
//   wr_ptr          rd_ptr
//   43210	      43210	(5-bit)
//   10000	      00000	(wr_ptr @ 16th location & rd_ptr @ 0th location)
//here, 4th bit of wr_ptr and 4th bit of rd_ptr are not equal and the rest of the bits are equal
assign full = ((wr_ptr[4] != rd_ptr[4]) && (wr_ptr[3:0] == rd_ptr[3:0]));

/*********************************************************************************************************************/

/*********************************************fifo lfd_state logic****************************************************/
/*reason for this delay will be explained in the top block*/

always@(posedge clock)
   begin
      if (!resetn)		//active low reset
         temp <= 0;
      else
         temp <= lfd_state;	//delaying lfd_state by 1 clock to latch the header byte
   end
   
/*********************************************************************************************************************/

/******************************************fifo write operation logic*************************************************/

always@(posedge clock)
   begin
      if (!resetn)			//active low reset
         begin
            for(i=0; i<16; i = i+1)
               mem[i] <= 0;		//all the memory locations of 9-bit wide should be made 0 for resetn = 0
               wr_ptr <= 0;		//write pointer points to the location 0
      	 end
      
      else if(soft_reset)		//active high soft reset - generated by SYNCHRONIZER block during the time out state of the ROUTER
         begin
            for(i=0; i<16; i = i+1)
               mem[i] <= 0;
               wr_ptr <= 0;
      	 end
      	 
      else if(write_enb && !full)	//if the fifo is not full and there is availability of some location and write_enb is enabled
         begin
            {mem[wr_ptr[3:0]][8], mem[wr_ptr[3:0]][7:0]} <= {temp, data_in};  //{wherever write pointer is pointing and 9th bit location(lfd_state bit), 
            									//wherever write pointer is pointing and 8 bit locations}
            wr_ptr <= wr_ptr + 1'b1;
         end
	end
       
/*********************************************************************************************************************/

/******************************************fifo internal counter logic************************************************/

always@(posedge clock)
   begin
      if(!resetn)
         count <= 0;
         
      else if(soft_reset)
         count <= 0;
         
      else if(mem[rd_ptr[3:0]][8] == 1)		//checking memory location that rd_ptr(4-bit) is pointing and 9th bit of this location is 1	(indication of Header byte)
         count <= mem[rd_ptr[3:0]][7:2] + 1'b1;	//internal counter loaded with Payload_length_of_packet + 1 (Parity byte)
         
      else if(read_enb && !empty)
         count <= count - 1'b1;
      else
         count <= count;
   end    
    
/*********************************************************************************************************************/

/*******************************************fifo read operation logic*************************************************/

always@(posedge clock)
   begin
      if(!resetn)
         begin
            data_out <= 0;
            rd_ptr <= 0;
         end
         
      else if(soft_reset)
            data_out <= 8'bz;
            
      else if(count == 0)				//which means Header + Payload + Parity are read
            data_out <= 8'bz;
                  
      else if(read_enb && !empty)
         begin
            data_out <= mem[rd_ptr[3:0]][7:0];	//memory w.r.t the rd_ptr that is pointing to [7:0] is sent as a data_out
            rd_ptr <= rd_ptr + 1'b1;
         end
      
      else
         data_out <= 8'bz;
   end
   
/*********************************************************************************************************************/

      
      
       
      
      
      
      
      
      
      
      
      
      
      
      
      
      
      
      
      
      



